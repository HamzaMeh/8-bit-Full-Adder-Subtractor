module tesben();
reg [3:0]a,b;
reg carry;
wire Cout;
reg [4:0]S;
wire [3:0]Y;

ALU alu(Cout,Y,a,b,carry,S);
initial begin
  //1
a[0]=0;a[1]=0;a[2]=0;a[3]=0;
b[0]=1;b[1]=0;b[2]=0;b[3]=0;
carry=0;
S[1]=0;S[0]=0;S[4]=0; 
#100 
//2
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
carry=1;
S[1]=0;S[0]=0;S[4]=0; 
#100 
//3
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[1]=0;S[0]=1;S[4]=0; 
#100 
//4
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[1]=1;S[0]=0;S[4]=0; 
#100 
//5
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[1]=1;S[0]=1;S[4]=0; 
#100
//6
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[2]=0;S[3]=0;S[4]=1; 
#100
//7
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[2]=1;S[3]=0;S[4]=1; 
#100 
//8
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[2]=0;S[3]=1;S[4]=1; 
#100 
//9
a[0]=0;a[1]=0;a[2]=1;a[3]=0;
b[0]=1;b[1]=1;b[2]=0;b[3]=0;
S[3]=1;S[2]=1;S[4]=1;  
end
endmodule